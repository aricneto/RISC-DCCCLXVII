module bindfiles;
    bind regfile_64 assert_type_r type_r (.*);
    bind instr_reg assert_type_r type_r (.*);
endmodule